// ECE:3350 SISC computer project
// Braden Miller & Scott Pearson

`timescale 1ns/100ps

module ctrl (clk, rst_f, opcode, mm, stat, rf_we, alu_op, wb_sel, pc_sel, pc_write, pc_rst, br_sel, ir_load);

  //I/O port declarations
  input clk, rst_f;
  input [3:0] opcode, mm, stat;
  output reg rf_we, wb_sel;
  output reg [3:0] alu_op;

  output reg pc_sel, pc_write, pc_rst; //pc control signals
  output reg br_sel; //br control signal
  output reg ir_load; //ir control signal

  
  // state parameter declarations
  
  parameter start0 = 0, start1 = 1, fetch = 2, decode = 3, execute = 4, mem = 5, writeback = 6;
   
  // opcode parameter declarations
  
  parameter NOOP = 0, REG_OP = 1, REG_IM = 2, SWAP = 3, BRA = 4, BRR = 5, BNE = 6, BNR = 7;
  parameter JPA = 8, JPR = 9, LOD = 10, STR = 11, CALL = 12, RET = 13, HLT = 15;
	
  // addressing modes
  
  parameter AM_IMM = 8;

  // state register and next state signal
  
  reg [2:0]  present_state, next_state;

  // initial procedure to initialize the present state to 'start0'.

  initial
    present_state = start0;

  /* Procedure that progresses the fsm to the next state on the positive edge of 
     the clock, OR resets the state to 'start1' on the negative edge of rst_f. 
     Notice that the computer is reset when rst_f is low, not high. */

  always @(posedge clk, negedge rst_f)
  begin
    if (rst_f == 1'b0)
      present_state <= start1;
    else
      present_state <= next_state;
  end
  
  /* The following combinational procedure determines the next state of the fsm. */

  always @(present_state, rst_f)
  begin
    case(present_state)
      start0:
        next_state = start1;
      start1:
	  if (rst_f == 1'b0) 
        next_state = start1;
	 else
         next_state = fetch;
      fetch:
        next_state = decode;
      decode:
        next_state = execute;
      execute:
        next_state = mem;
      mem:
        next_state = writeback;
      writeback:
        next_state = fetch;
      default:
        next_state = start1;
    endcase
  end

  //Update control signal outputs depending on state and opcode
  always @(present_state, opcode, mm) //got rid of stat
  begin

  // Default value of 0 for output control signals
  rf_we = 1'b0;
  alu_op = 4'b0000;
  wb_sel = 1'b0;

  pc_sel = 1'b0;   //pc_sel = 1 increments program counter
  pc_write = 1'b0; //pc_write: When this control bit changes to 1, the selected value (either
          		 //the branch address or PC+1) is saved to pc_out and held there until
          		 //the next time pc_en is set to 1.
  pc_rst = 1'b0;   //resets program counter
  br_sel = 1'b0;   //(relative branch, br_sel = 0) or to add it to 0 (absolute branch, br_sel = 1).
  ir_load = 1'b0;  //ir_load: if ir_load is = 1, the IR is loaded with read_data
  
  case(present_state)
        start1: 
        begin
          pc_rst = 1'b1;   // Reset PC when in start1 state
   	end
    
    fetch:
    begin
      ir_load = 1'b1;  // Load instruction register in fetch state
   //may not need   pc_sel = 1'b0;   // Select PC+1
      pc_write = 1'b1; // Update PC with PC+1
    end


      decode:
      begin
        // Determine branch selection and PC write based on branch instructions
        case(opcode)
          BRA, JPA, CALL: begin
            pc_sel = 1'b1;  // Select branch address
            br_sel = 1'b1;  // Absolute branch/jump
            if (opcode == BRA) begin
              // Branch if mm & stat is not zero
              pc_write = ((mm & stat) != 4'b0000);
            end
            else begin
              // Always jump for JPA and CALL
              pc_write = 1'b1;
            end
          end

          BRR, JPR, RET: begin
            pc_sel = 1'b1;  // Select branch address
            br_sel = 1'b0;  // Relative branch
            if (opcode == BRR) begin
              // Branch if mm & stat is not zero
              pc_write = ((mm & stat) != 4'b0000);
            end
            else begin
              // Always jump for JPR and RET
              pc_write = 1'b1;
            end
          end

          BNE: begin
            pc_sel = 1'b1;   // Select branch address
            br_sel = 1'b1;   // Absolute branch
            // Write PC if condition is met (mm & stat is zero)
            pc_write = ((mm & stat) == 4'b0000);
          end

          BNR: begin
            pc_sel = 1'b1;   // Select branch address
            br_sel = 1'b0;   // Relative branch
            // Write PC if condition is met (mm & stat is zero)
            pc_write = ((mm & stat) == 4'b0000);
          end
        endcase
      end
	

	execute:
	begin
	 if(opcode == REG_OP)
	    alu_op = 4'b0001; //if opcode is reg_op, set alu_op to 0001
	 if(opcode == REG_IM)
	    alu_op = 4'b0011; //if opcode is reg_im, set alu_op to 0011
	end

	mem:
	begin
	 if(opcode == REG_OP)
	    alu_op = 4'b0000; //if opcode is reg_op, set alu_op to 0000
	 if(opcode == REG_IM)
	    alu_op = 4'b0010; //if opcode is reg_im, set alu_op to 0010
	end

	writeback:
	begin
	   if (opcode == REG_OP || opcode == REG_IM)
		rf_we = 1'b1; //set rf_we to 1 if opcode is REG_OP or REG_IM
	end

	default: 
	begin
	 rf_we = 1'b0; //reset re_we back to default
	 wb_sel = 1'b0;
         alu_op = 4'b0000;
         pc_sel = 1'b0;
         pc_write = 1'b0;
         pc_rst = 1'b0;
         br_sel = 1'b0;
         ir_load = 1'b0;
	end
     endcase
  end

    



// Halt on HLT instruction
  always @ (opcode)
  begin
    if (opcode == HLT)
    begin 
      #5 $display ("Halt."); //Delay 5 ns so $monitor will print the halt instruction
      $stop;
    end
  end
    
  
endmodule
